module Mod2(input clk,
    input  io_in02,
    output io_out02
);



  assign io_out02 = io_in02;
endmodule
