module prova01(
    input  io_A,
    output io_B
);



  assign io_B = io_A;
endmodule

